library verilog;
use verilog.vl_types.all;
entity maq_refri_tb is
end maq_refri_tb;
